library verilog;
use verilog.vl_types.all;
entity tb_rightshifter is
end tb_rightshifter;
