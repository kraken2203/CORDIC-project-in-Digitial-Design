library verilog;
use verilog.vl_types.all;
entity tb_stage0 is
end tb_stage0;
